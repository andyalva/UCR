module test
(output f,
input a, b);
and A(f, a, b);
endmodule